interface intf(input clk);
  reg reset;
  reg [2:0] d;
  reg [2:0]q;
endinterface
